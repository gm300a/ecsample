module pllcut(input clk,rst,a,output clko,x) ;
    
